`ifdef VEDIT
  `include "vedit_inc.v"
`endif
